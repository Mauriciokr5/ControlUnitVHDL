LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALU IS

	PORT (
		  ENTRADA:IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		  ENTRADAB: IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		  SEL4:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  OUT_ALU:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		  SIGNO,INDET:OUT STD_LOGIC)
		  ;
			
END ALU;

ARCHITECTURE ALUB OF ALU IS
	
	SIGNAL SEL:STD_LOGIC_VECTOR(1 DOWNTO 0):="00";--SELEC DEL MUX;
	SIGNAL NBIN: STD_LOGIC_VECTOR(13 DOWNTO 0):="00000000000000";
	SIGNAL NBIN_AUX: STD_LOGIC_VECTOR(13 DOWNTO 0):="00000000000000";--NUMERO BINARIO 14 BITS
	SIGNAL S_B:STD_LOGIC_VECTOR(11 DOWNTO 0):="000000000000";--SE�AL PARA ALAMCENAR A "B"
	SIGNAL S_BAUX:STD_LOGIC_VECTOR(12 DOWNTO 0);--SE�AL QUE SE ENVIARA AL SUMADOR DE 13 BITS
	SIGNAL S_A:STD_LOGIC_VECTOR(11 DOWNTO 0):="000000000000";--SE�AL PARA ALAMCENAR A "A"
	SIGNAL S_AAUX:STD_LOGIC_VECTOR(12 DOWNTO 0);--SE�AL QUE SE ENVIARA AL SUMADOR DE 13 BITS
	SIGNAL RESTA8:STD_LOGIC;
	SIGNAL RESTA12:STD_LOGIC;
	SIGNAL FACT1: STD_LOGIC_VECTOR(5 DOWNTO 0); --SE ENVIA AL MUL.
	SIGNAL FACT2:STD_LOGIC_VECTOR(5 DOWNTO 0);-- ENVIAR AL  MUL.
	SIGNAL RESULT:STD_LOGIC_VECTOR(11 DOWNTO 0):="000000000000";--N B 12B
	SIGNAL COCIENTE:STD_LOGIC_VECTOR (5 DOWNTO 0);
	SIGNAL DIV:STD_LOGIC;
	SIGNAL LED_AUX:STD_LOGIC_VECTOR(12 DOWNTO 0);
	SIGNAL S_INDET:STD_LOGIC;
	SIGNAL BCDAUX: STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL temp_LED_AUX:STD_LOGIC_VECTOR(12 DOWNTO 0);
	COMPONENT SUMADOR_13BITS IS

	PORT(A,B:IN STD_LOGIC_VECTOR(12 DOWNTO 0);
		 S:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		 COUT12:OUT STD_LOGIC);
		
	END COMPONENT;
	
	COMPONENT mult_comb_gen is
	Generic ( g_bits : natural := 6 ); 
	Port (fact1 : in STD_LOGIC_VECTOR (g_bits-1 downto 0); 
		  fact2 : in STD_LOGIC_VECTOR (g_bits-1 downto 0); 
		  prod : out STD_LOGIC_VECTOR (2*g_bits-1 downto 0)); -- doble de bits para el producto
	end COMPONENT;
	
	COMPONENT BRRL_S IS 
	PORT(SEL:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 PIN:IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 POUT:OUT STD_LOGIC_VECTOR(12 DOWNTO 0)); 
	END COMPONENT;
	
	COMPONENT DIV6 IS 
	PORT(DIVIDENDO,DIVISOR:IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 COCIENTE:OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		 INDET: OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT convertidor_BCD is 
	PORT(
	bin: in std_logic_vector(12 downto 0);
	bcd: out std_logic_vector(15 downto 0)
	);
	end COMPONENT;
	
	COMPONENT display_4digitos is
	port(
		CLK: in std_logic;
		in_bcd: in std_logic_vector(15 downto 0);
		sel_d: out std_logic_vector(3 downto 0);
		seg_d: out std_logic_vector(6 downto 0)
		);
	end COMPONENT;

	
BEGIN 
	
	--AQUI SE HACE LA SELECCION DE OPERACION
	OPERACION:PROCESS (SEL4,ENTRADA, ENTRADAB,RESTA8,RESTA12)
		BEGIN
			S_A<=ENTRADA;
			S_B <= ENTRADAB;
			RESTA8<='0';
			RESTA12<='0';
			CASE SEL4 IS
				-- COMPLEMENTO A 1 DE A
				WHEN "0001" => temp_LED_AUX <= '0' & NOT(S_A); 
				-- COMPLEMENTO A 2 DE A
				WHEN "0010" => temp_LED_AUX <= (NOT('0' & S_A)+'1');
				-- AND ENTRE A Y B
				WHEN "0011" => temp_LED_AUX <= '0' & (S_A AND S_B);
				-- OR ENTRE A Y B
				WHEN "0100" => temp_LED_AUX <= '0' & (S_A OR S_B);
				-- LSL
				WHEN "0101" => temp_LED_AUX <=LED_AUX;
				-- SUMA DE 1 BYTE C/ CARRY OUT
				WHEN "0111" => S_AAUX <= "00000"& S_A(7 DOWNTO 0);
							   S_BAUX <= "00000"& S_B(7 DOWNTO 0);
				-- RESTA DE 1 BYTE C/ CARRY OUT
				WHEN "1000" => S_AAUX <= "00000"& ENTRADA(7 DOWNTO 0);
								S_BAUX <= ("11111" & NOT S_B(7 DOWNTO 0))+'1';
								RESTA8<='1';
				--MULTIPLICACION 5 BITS
				WHEN "1001" => FACT1<=ENTRADA(5 DOWNTO 0); -- A*B(6 BITS)
								FACT2 <= ENTRADAB(5 DOWNTO 0);
								--S_AAUX<= '0' & RESULT;
								--S_BAUX<="0000000000000";
				--DIVISION 5 BITS		
				WHEN "1010" => S_AAUX <= "0000000" & COCIENTE ;-- A/B(6 BITS)	
								S_BAUX <= "0000000000000";
								DIV<='1';
								
				WHEN OTHERS => temp_LED_AUX<=LED_AUX; --CORRIMIRENTO IZQ.	

			END CASE;
	END PROCESS OPERACION;
	
	CALL1: BRRL_S PORT MAP (SEL=>S_B(3 DOWNTO 0),PIN=>S_A,POUT=>LED_AUX);
	--COMPONENTE MULTIPLICADOR
	CALL2:mult_comb_gen GENERIC MAP(G_BITS=>6)PORT MAP(fact1=>fact1,fact2=>fact2,prod=>RESULT);	 
	--DIVISOR
	CALL4: DIV6 PORT MAP(DIVIDENDO=>S_A(5 DOWNTO 0),DIVISOR=>S_B(5DOWNTO 0),COCIENTE=>COCIENTE,INDET=>S_INDET); 
		-- PORT MAP DEL SUMADOR 13 BITS
	CALL0: SUMADOR_13BITS PORT MAP(A=>S_AAUX,B=>S_BAUX,S=>NBIN_AUX(12 DOWNTO 0),COUT12=>NBIN_AUX(13));
	 
	OUT_ALU <= '0' & RESULT;
END ALUB;