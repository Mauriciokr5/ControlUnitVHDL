LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUMADOR_COMPLETO IS

	PORT(A,B,CIN:IN STD_LOGIC;
		 S,COUT:OUT STD_LOGIC);
		 
END ENTITY;

ARCHITECTURE COMPORTAMIENTO OF SUMADOR_COMPLETO IS
	
	SIGNAL S_XOR:STD_LOGIC;
	SIGNAL S_AND1:STD_LOGIC;
	SIGNAL S_AND2:STD_LOGIC;
	SIGNAL S_OR:STD_LOGIC;

BEGIN

	S_XOR <= A XOR B;
	S_AND1<= A AND B;
	S_OR <= A OR B;
	S_AND2 <=S_OR AND CIN;
	S <= S_XOR XOR CIN;
	COUT <= S_AND1 OR S_AND2;
	
END ARCHITECTURE;
