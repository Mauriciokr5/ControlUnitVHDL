LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUMADOR_13BITS IS

	PORT(A,B:IN STD_LOGIC_VECTOR(12 DOWNTO 0);
		 S:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		 COUT12:OUT STD_LOGIC);
		
END ENTITY;

ARCHITECTURE COMPORTAMIENTO OF SUMADOR_13BITS IS

	COMPONENT SUMADOR_COMPLETO IS

		PORT(A,B,CIN:IN STD_LOGIC;
			S,COUT:OUT STD_LOGIC);

		END COMPONENT;

	SIGNAL COUT0,COUT1,COUT2:STD_LOGIC;
	SIGNAL COUT3,COUT4,COUT5:STD_LOGIC;
	SIGNAL COUT6,COUT7,COUT8:STD_LOGIC;
	SIGNAL COUT9,COUT10,COUT11:STD_LOGIC;
	
BEGIN

LLAMADA0:SUMADOR_COMPLETO PORT MAP (A=>A(0),B=>B(0),CIN=>'0',S=>S(0),COUT=>COUT0);
LLAMADA1:SUMADOR_COMPLETO PORT MAP (A=>A(1),B=>B(1),CIN=>COUT0,S=>S(1),COUT=>COUT1);
LLAMADA2:SUMADOR_COMPLETO PORT MAP (A=>A(2),B=>B(2),CIN=>COUT1,S=>S(2),COUT=>COUT2);
LLAMADA3:SUMADOR_COMPLETO PORT MAP (A=>A(3),B=>B(3),CIN=>COUT2,S=>S(3),COUT=>COUT3);
LLAMADA4:SUMADOR_COMPLETO PORT MAP (A=>A(4),B=>B(4),CIN=>COUT3,S=>S(4),COUT=>COUT4);
LLAMADA5:SUMADOR_COMPLETO PORT MAP (A=>A(5),B=>B(5),CIN=>COUT4,S=>S(5),COUT=>COUT5);
LLAMADA6:SUMADOR_COMPLETO PORT MAP (A=>A(6),B=>B(6),CIN=>COUT5,S=>S(6),COUT=>COUT6);
LLAMADA7:SUMADOR_COMPLETO PORT MAP (A=>A(7),B=>B(7),CIN=>COUT6,S=>S(7),COUT=>COUT7);
LLAMADA8:SUMADOR_COMPLETO PORT MAP (A=>A(8),B=>B(8),CIN=>COUT7,S=>S(8),COUT=>COUT8);
LLAMADA9:SUMADOR_COMPLETO PORT MAP (A=>A(9),B=>B(9),CIN=>COUT8,S=>S(9),COUT=>COUT9);
LLAMADA10:SUMADOR_COMPLETO PORT MAP (A=>A(10),B=>B(10),CIN=>COUT9,S=>S(10),COUT=>COUT10);
LLAMADA11:SUMADOR_COMPLETO PORT MAP (A=>A(11),B=>B(11),CIN=>COUT9,S=>S(11),COUT=>COUT11);
LLAMADA12:SUMADOR_COMPLETO PORT MAP (A=>A(12),B=>B(12),CIN=>COUT10,S=>S(12),COUT=>COUT12);

END ARCHITECTURE;