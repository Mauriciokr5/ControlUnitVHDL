LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY BRRL_S IS 
	PORT(SEL:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 PIN:IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 POUT:OUT STD_LOGIC_VECTOR(12 DOWNTO 0)); 
END BRRL_S;

ARCHITECTURE BRRL_S_B OF BRRL_S IS
	BEGIN
		PROCESS (SEL,PIN)
		BEGIN
 
		CASE SEL IS 

			WHEN "0000" => POUT <= '0' & PIN; --NECESARIO PARA CORRIMIENTO 0
			WHEN "0001" => POUT <= '0' & PIN(10 DOWNTO 0) & '0';
			WHEN "0010" => POUT <= '0' & PIN(9 DOWNTO 0) & "00";
			WHEN "0011" => POUT <= '0' & PIN(8 DOWNTO 0) & "000";
			WHEN "0100" => POUT <= '0' & PIN(7 DOWNTO 0) & "0000";
			WHEN "0101" => POUT <= '0' & PIN(6 DOWNTO 0) & "00000";
			WHEN "0110" => POUT <= '0' & PIN(5 DOWNTO 0) & "000000";
			WHEN "0111" => POUT <= '0' & PIN(4 DOWNTO 0) & "0000000";
			WHEN "1000" => POUT <= '0' & PIN(3 DOWNTO 0) & "00000000";
			WHEN "1001" => POUT <= '0' & PIN(2 DOWNTO 0) & "000000000";
			WHEN "1010" => POUT <= '0' & PIN(1 DOWNTO 0) &"0000000000";
			WHEN "1011" => POUT <= '0' & PIN(0) & "00000000000";
			WHEN OTHERS => POUT<= "0000000000000";
		END CASE;
		END PROCESS;
END BRRL_S_B;